
module buffer(A,O);
input A;
output O;
buf bu(O,A);
endmodule
